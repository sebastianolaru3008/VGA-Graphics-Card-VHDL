library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity image_graph is
	port(
		img_e: in std_logic;
		pixel_x, pixel_y: in std_logic_vector(9 downto 0);
		c_sel: in std_logic_vector(1 downto 0);
		p_sel: in std_logic_vector(1 downto 0);
		rgb:  out std_logic_vector(7 downto 0) 	
		);
end image_graph;

architecture behave of image_graph is 

signal pix_x, pix_y: unsigned(9 downto 0);
constant MAX_X : integer := 640;  
constant MAX_Y : integer := 480;
constant SPRITE_SIZE: integer:= 64;	

constant sprite_x_l: unsigned(9 downto 0) := to_unsigned(MAX_X-SPRITE_SIZE-1,10);
constant sprite_x_r: unsigned(9 downto 0) := to_unsigned(MAX_X-1,10); 
constant sprite_y_t: unsigned(9 downto 0) := to_unsigned(MAX_Y-SPRITE_SIZE-1,10);
constant sprite_y_b: unsigned(9 downto 0) := to_unsigned(MAX_Y-1,10);

type rom_type is array(0 to 63) of std_logic_vector(0 to 63);
signal rom_row, rom_col: unsigned(5 downto 0);
signal rom_data: std_logic_vector(63 downto 0);
signal rom_bit: std_logic;
signal rb_sprite_on, inside_sprite_on: std_logic;
																  
constant HEART: rom_type:= (									  
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000001111111110000000000000000000000111111111000000000000",
"0000000000111111111111100000000000000000011111111111110000000000",
"0000000011111111111111111000000000000001111111111111111100000000",
"0000001111111111111111111110000000000111111111111111111111000000",
"0000011111111111111111111111000000001111111111111111111111100000",
"0000111111111111111111111111100000011111111111111111111111110000",
"0001111111111111111111111111110000111111111111111111111111111000",
"0001111111111111111111111111110000111111111111111111111111111000",
"0011111111111111111111111111111001111111111111111111111111111100",
"0011111111111111111111111111111001111111111111111111111111111100",
"0111111111111111111111111111111111111111111111111111111111111110",
"0111111111111111111111111111111111111111111111111111111111111110",
"1111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111",
"0111111111111111111111111111111111111111111111111111111111111110",
"0111111111111111111111111111111111111111111111111111111111111110",
"0011111111111111111111111111111111111111111111111111111111111100",
"0011111111111111111111111111111111111111111111111111111111111100",
"0001111111111111111111111111111111111111111111111111111111111000",
"0001111111111111111111111111111111111111111111111111111111111000",
"0000111111111111111111111111111111111111111111111111111111110000",
"0000011111111111111111111111111111111111111111111111111111100000",
"0000001111111111111111111111111111111111111111111111111111000000",
"0000000111111111111111111111111111111111111111111111111110000000",
"0000000011111111111111111111111111111111111111111111111100000000",
"0000000001111111111111111111111111111111111111111111111000000000",
"0000000000111111111111111111111111111111111111111111110000000000",
"0000000000011111111111111111111111111111111111111111100000000000",
"0000000000001111111111111111111111111111111111111111000000000000",
"0000000000000111111111111111111111111111111111111110000000000000",
"0000000000000011111111111111111111111111111111111100000000000000",
"0000000000000001111111111111111111111111111111111000000000000000",
"0000000000000000111111111111111111111111111111110000000000000000",
"0000000000000000011111111111111111111111111111100000000000000000",
"0000000000000000001111111111111111111111111111000000000000000000",
"0000000000000000000111111111111111111111111110000000000000000000",
"0000000000000000000011111111111111111111111100000000000000000000",
"0000000000000000000001111111111111111111111000000000000000000000",
"0000000000000000000000111111111111111111110000000000000000000000",
"0000000000000000000000011111111111111111100000000000000000000000",
"0000000000000000000000001111111111111111000000000000000000000000",
"0000000000000000000000000111111111111110000000000000000000000000",
"0000000000000000000000000011111111111100000000000000000000000000",
"0000000000000000000000000001111111111000000000000000000000000000",
"0000000000000000000000000000111111110000000000000000000000000000",
"0000000000000000000000000000011111100000000000000000000000000000",
"0000000000000000000000000000001111000000000000000000000000000000",
"0000000000000000000000000000000110000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000");
																  
constant CHERIES: rom_type:= (										  
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000001111111111110000000000000000000000",
"0000000000000000000000000000001111111111110000000000000000000000",
"0000000000000000000000000000001111111111110000000000000000000000",
"0000000000000000000000000000011111111111110000000000000000000000",
"0000000000000000000000000001100000100000000000000000000000000000",
"0000000000000000000000000001000001000000000000000000000000000000",
"0000000000000000000000000001000001000000000000000000000000000000",
"0000000000000000000000000010000001000000000000000000000000000000",
"0000000000000000000000000010000001000000000000000000000000000000",
"0000000000000000000000000100000001000000000000000000000000000000",
"0000000000000000000000000100000000100000000000000000000000000000",
"0000000000000000000000000100000000100000000000000000000000000000",
"0000000000000000000000000100000000100000000000000000000000000000",
"0000000000000000000000001000000000010000000000000000000000000000",
"0000000000000000000000001000000000001000000000000000000000000000",
"0000000000000000000000001000000000001100000000000000000000000000",
"0000000000000000000000010000000000000010000000000000000000000000",
"0000000000000000000000010000000000000011000000000000000000000000",
"0000000000000000000000010000000000000001100000000000000000000000",
"0000000000000000000000010000000000000000110000000000000000000000",
"0000000000000000000000111000000000000000011100000000000000000000",
"0000000000000000000000111000000000000000011100000000000000000000",
"0000000000000000000011111110000000000001111111000000000000000000",
"0000000000000000001111111111100000000111111111110000000000000000",
"0000000000000000011111111111110000001111111111111000000000000000",
"0000000000000000111111111111111000011111111111111100000000000000",
"0000000000000001111111111111111100111111111111111110000000000000",
"0000000000000001111111111111111100111111111111111110000000000000",
"0000000000000011111111111111111111111111111111111111000000000000",
"0000000000000011111111111111111111111111111111111111000000000000",
"0000000000000011111111111111111111111111111111111111000000000000",
"0000000000000011111111111111111111111111111111111111000000000000",
"0000000000000011111111111111111111111111111111111111000000000000",
"0000000000000011111111111111111111111111111111111111000000000000",
"0000000000000011111111111111111111111111111111111111000000000000",
"0000000000000001111111111111111100111111111111111110000000000000",
"0000000000000001111111111111111100111111111111111110000000000000",
"0000000000000000111111111111111000011111111111111100000000000000",
"0000000000000000011111111111110000001111111111111000000000000000",
"0000000000000000001111111111100000000111111111110000000000000000",
"0000000000000000000011111110000000000001111111000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000");

constant BALL: rom_type:= (
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000001111111111100000000000000000000000000",
"0000000000000000000000001111111111111111100000000000000000000000",
"0000000000000000000001111111111111111111111100000000000000000000",
"0000000000000000000111111111111111111111111111000000000000000000",
"0000000000000000001111111111111111111111111111100000000000000000",
"0000000000000000111111111111111111111111111111111000000000000000",
"0000000000000001111111111111111111111111111111111100000000000000",
"0000000000000011111111111111111111111111111111111110000000000000",
"0000000000000111111111111111111111111111111111111111000000000000",
"0000000000001111111111111111111111111111111111111111100000000000",
"0000000000011111111111111111111111111111111111111111110000000000",
"0000000000111111111111111111111111111111111111111111111000000000",
"0000000000111111111111111111111111111111111111111111111000000000",
"0000000001111111111111111111111111111111111111111111111100000000",
"0000000011111111111111111111111111111111111111111111111110000000",
"0000000011111111111111111111111111111111111111111111111110000000",
"0000000111111111111111111111111111111111111111111111111111000000",
"0000000111111111111111111111111111111111111111111111111111000000",
"0000000111111111111111111111111111111111111111111111111111000000",
"0000001111111111111111111111111111111111111111111111111111100000",
"0000001111111111111111111111111111111111111111111111111111100000",
"0000001111111111111111111111111111111111111111111111111111100000",
"0000011111111111111111111111111111111111111111111111111111110000",
"0000011111111111111111111111111111111111111111111111111111110000",
"0000011111111111111111111111111111111111111111111111111111110000",
"0000011111111111111111111111111111111111111111111111111111110000",
"0000011111111111111111111111111111111111111111111111111111110000",
"0000011111111111111111111111111111111111111111111111111111110000",
"0000011111111111111111111111111111111111111111111111111111110000",
"0000011111111111111111111111111111111111111111111111111111110000",
"0000011111111111111111111111111111111111111111111111111111110000",
"0000011111111111111111111111111111111111111111111111111111110000",
"0000011111111111111111111111111111111111111111111111111111110000",
"0000001111111111111111111111111111111111111111111111111111100000",
"0000001111111111111111111111111111111111111111111111111111100000",
"0000001111111111111111111111111111111111111111111111111111100000",
"0000000111111111111111111111111111111111111111111111111111000000",
"0000000111111111111111111111111111111111111111111111111111000000",
"0000000111111111111111111111111111111111111111111111111111000000",
"0000000011111111111111111111111111111111111111111111111110000000",
"0000000011111111111111111111111111111111111111111111111110000000",
"0000000001111111111111111111111111111111111111111111111100000000",
"0000000000111111111111111111111111111111111111111111111000000000",
"0000000000111111111111111111111111111111111111111111111000000000",
"0000000000011111111111111111111111111111111111111111110000000000",
"0000000000001111111111111111111111111111111111111111100000000000",
"0000000000000111111111111111111111111111111111111111000000000000",
"0000000000000011111111111111111111111111111111111110000000000000",
"0000000000000001111111111111111111111111111111111100000000000000",
"0000000000000000111111111111111111111111111111111000000000000000",
"0000000000000000001111111111111111111111111111100000000000000000",
"0000000000000000000111111111111111111111111111000000000000000000",
"0000000000000000000001111111111111111111111100000000000000000000",
"0000000000000000000000001111111111111111100000000000000000000000",
"0000000000000000000000000001111111111100000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000");
																  
constant INVADER: rom_type:= (								 
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000011111100000000000000000000000000000011111100000000000",
"0000000000011111100000000000000000000000000000011111100000000000",
"0000000000011111100000000000000000000000000000011111100000000000",
"0000000000011111100000000000000000000000000000011111100000000000",
"0000000000011111100000000000000000000000000000011111100000000000",
"0000000000011111100000000000000000000000000000011111100000000000",
"0000000000000000011111100000000000000000011111100000000000000000",
"0000000000000000011111100000000000000000011111100000000000000000",
"0000000000000000011111100000000000000000011111100000000000000000",
"0000000000000000011111100000000000000000011111100000000000000000",
"0000000000000000011111100000000000000000011111100000000000000000",
"0000000000000000011111100000000000000000011111100000000000000000",
"0000000000011111111111111111111111111111111111111111100000000000",
"0000000000011111111111111111111111111111111111111111100000000000",
"0000000000011111111111111111111111111111111111111111100000000000",
"0000000000011111111111111111111111111111111111111111100000000000",
"0000000000011111111111111111111111111111111111111111100000000000",
"0000000000011111111111111111111111111111111111111111100000000000",
"0000011111111111100000011111111111111111100000011111111111100000",
"0000011111111111100000011111111111111111100000011111111111100000",
"0000011111111111100000011111111111111111100000011111111111100000",
"0000011111111111100000011111111111111111100000011111111111100000",
"0000011111111111100000011111111111111111100000011111111111100000",
"0000011111111111100000011111111111111111100000011111111111100000",
"1111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111",
"1111100000011111111111111111111111111111111111111111100000011111",
"1111100000011111111111111111111111111111111111111111100000011111",
"1111100000011111111111111111111111111111111111111111100000011111",
"1111100000011111111111111111111111111111111111111111100000011111",
"1111100000011111111111111111111111111111111111111111100000011111",
"1111100000011111111111111111111111111111111111111111100000011111",
"1111100000011111100000000000000000000000000000011111100000011111",
"1111100000011111100000000000000000000000000000011111100000011111",
"1111100000011111100000000000000000000000000000011111100000011111",
"1111100000011111100000000000000000000000000000011111100000011111",
"1111100000011111100000000000000000000000000000011111100000011111",
"1111100000011111100000000000000000000000000000011111100000011111",
"0000000000000000011111111111100000011111111111100000000000000000",
"0000000000000000011111111111100000011111111111100000000000000000",
"0000000000000000011111111111100000011111111111100000000000000000",
"0000000000000000011111111111100000011111111111100000000000000000",
"0000000000000000011111111111100000011111111111100000000000000000",
"0000000000000000011111111111100000011111111111100000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000");
																  
		   														  
begin  	 
	pix_x <= unsigned(pixel_x);
	pix_y <= unsigned(pixel_y);	 
	
	process	(pix_x,pix_y)
	begin
		if (sprite_x_l <= pix_x) and (pix_x <= sprite_x_r) and (sprite_y_t <= pix_y) and (pix_y <= sprite_y_b) then
			inside_sprite_on <= '1';
		else 
			inside_sprite_on <= '0'; 
		end if;
	end process;
	
	rom_row <= pix_y(5 downto 0) - sprite_y_t(5 downto 0); -- because they are close in vlaue if inside is true	 
	rom_col <= pix_x(5 downto 0) - sprite_x_l(5 downto 0); -- same here
	
	
	rom_data <= HEART(to_integer(rom_row))   when p_sel = "00"
	else CHERIES(to_integer(rom_row)) when p_sel = "01"
	else BALL(to_integer(rom_row)) when p_sel = "10"  
	else INVADER(to_integer(rom_row)); 
		
	rom_bit <= rom_data(to_integer(rom_col));
	rb_sprite_on <= '1' when (inside_sprite_on = '1') and (rom_bit = '1') else '0';
					  
		
	process (img_e, c_sel, rb_sprite_on)
		begin
			if(img_e = '1' and rb_sprite_on = '1') then
				if   (c_sel = "00") then rgb <= "11111111";
				elsif(c_sel = "01") then rgb <= "11111100";
				elsif(c_sel = "10") then rgb <= "00000011";
				elsif(c_sel = "11") then rgb <= "11100011";
				end if;
			else
				rgb <= "00000000";
			end if;
	end process;
	
end architecture;